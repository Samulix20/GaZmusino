/* verilator lint_off UNUSEDSIGNAL */

module testbench (
    input logic clk, resetn
);


endmodule
